`include "config.v"

module mem_ctrl (
    input  wire clk,
    input  wire rst,
    input  wire rdy,

    //ram
    input  wire ram_din,
    output reg 
);

endmodule //mem_ctrl